/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  // assign uio_out = 0;
  // assign uio_oe  = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};
    wire more_unused = &{ui_in, uio_in};

    // 3-bit counter with tristate output
    reg [2:0] count;
    
    // Synchronous counter logic with reset
    always @(posedge clk) begin
        if (!rst_n)
            // Reset to 0 if press reset
            count <= 3'b000;
        else
            count <= count + 1;
    end
    
    // Tristate output buffer, let ui_in[0] be the enable signal
    assign temp = {5'b00000, count};
    assign uo_out = ui_in[0] ? temp : '8bz
    assign uio_out = 0;
    assign uio_oe = 0;

endmodule
